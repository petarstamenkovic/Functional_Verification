library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity rom is
    generic (WIDTH: positive := 32;
             SIZE: positive := 180;
			 SIZE_WIDTH: positive := 8);
    port (clk_a : in std_logic;
          clk_b : in std_logic;
          en_a: in std_logic;
          en_b: in std_logic;
          addr_a : in std_logic_vector(SIZE_WIDTH - 1 downto 0);
          addr_b : in std_logic_vector(SIZE_WIDTH - 1 downto 0);
          data_a_o: out std_logic_vector(WIDTH - 1 downto 0);
          data_b_o: out std_logic_vector(WIDTH - 1 downto 0));
end rom;

architecture Behavioral of rom is
    type rom_type is array(0 to SIZE - 1) of std_logic_vector(WIDTH - 1 downto 0);
    signal ROM : rom_type := (
            "00000000000000000100000000000000", "00000001000111010011111111111101", "00000010001110110011111111110110", "00000011010110010011111111101001", 
			"00000100011101100011111111011000", "00000101100100110011111111000001", "00000110101100000011111110100110", "00000111110011000011111110000101", 
			"00001000111010000011111101100000", "00001010000000110011111100110110", "00001011000111010011111100000111", "00001100001101100011111011010010", 
			"00001101010011100011111010011001", "00001110011001010011111001011100", "00001111011110110011111000011001", "00010000100100000011110111010001", 
			"00010001101001000011110110000101", "00010010101101100011110100110100", "00010011110001100011110011011110", "00010100110101100011110010000011", 
			"00010101111000110011110000100011", "00010110111011110011101110111111", "00010111111110010011101101010110", "00011001000000010011101011101001", 
			"00011010000001110011101001110111", "00011011000011000011101000000000", "00011100000011100011100110000101", "00011101000011100011100100000110", 
			"00011110000010110011100010000010", "00011111000001110011011111111001", "00011111111111110011011101101100", "00100000111101100011011011011011", 
			"00100001111010100011011001000110", "00100010110110110011010110101100", "00100011110010010011010100001110", "00100100101101010011010001101100", 
			"00100101100111100011001111000110", "00100110100001000011001100011100", "00100111011001100011001001101110", "00101000010001100011000110111100", 
			"00101001001000110011000100000110", "00101001111111000011000001001101", "00101010110100110010111110001111", "00101011101001010010111011001110", 
			"00101100011101010010111000001001", "00101101010000010010110101000001", "00101110000010010010110001110101", "00101110110011100010101110100101", 
			"00101111100011110010101011010011", "00110000010011010010100111111100", "00110001000001100010100100100011", "00110001101111000010100001000110", 
			"00110010011011100010011101100110", "00110011000111000010011010000100", "00110011110001100010010110011110", "00110100011011000010010010110101", 
			"00110101000011100010001111001001", "00110101101011000010001011011011", "00110110010001100010000111101010", "00110110110110110010000011110110", 
			"00110111011011000010000000000000", "00110111111110010001111100000111", "00111000100000100001111000001011", "00111001000001100001110100001110", 
			"00111001100001010001110000001110", "00111010000000000001101100001100", "00111010011101110001101000000111", "00111010111010010001100100000001", 
			"00111011010101100001011111111001", "00111011101111110001011011101111", "00111100001000110001010111100011", "00111100100000110001010011010110", 
			"00111100110111100001001111000110", "00111101001101000001001010110110", "00111101100001010001000110100100", "00111101110100010001000010010000", 
			"00111110000110010000111101111011", "00111110010111000000111001100101", "00111110100110010000110101001110", "00111110110100100000110000110110", 
			"00111111000001110000101100011101", "00111111001101100000101000000011", "00111111011000000000100011101000", "00111111100001010000011111001100", 
			"00111111101001100000011010110000", "00111111110000010000010110010011", "00111111110110000000010001110110", "00111111111010010000001101011001", 
			"00111111111101100000001000111011", "00111111111111010000000100011101", "01000000000000000000000000000000", "00111111111111011111111011100010", 
			"00111111111101101111110111000100", "00111111111010011111110010100110", "00111111110110001111101110001001", "00111111110000011111101001101100", 
			"00111111101001101111100101001111", "00111111100001011111100000110011", "00111111011000001111011100010111", "00111111001101101111010111111100", 
			"00111111000001111111010011100010", "00111110110100101111001111001001", "00111110100110011111001010110001", "00111110010111001111000110011010", 
			"00111110000110011111000010000100", "00111101110100011110111101101111", "00111101100001011110111001011011", "00111101001101001110110101001001", 
			"00111100110111101110110000111001", "00111100100000111110101100101001", "00111100001000111110101000011100", "00111011101111111110100100010000", 
			"00111011010101101110100000000110", "00111010111010011110011011111110", "00111010011101111110010111111000", "00111010000000001110010011110011", 
			"00111001100001011110001111110001", "00111001000001101110001011110001", "00111000100000101110000111110100", "00110111111110011110000011111000", 
			"00110111011011001110000000000000", "00110110110110111101111100001001", "00110110010001101101111000010101", "00110101101011001101110100100100", 
			"00110101000011101101110000110110", "00110100011011001101101101001010", "00110011110001101101101001100001", "00110011000111001101100101111011", 
			"00110010011011101101100010011001", "00110001101111001101011110111001", "00110001000001101101011011011100", "00110000010011011101011000000011", 
			"00101111100011111101010100101100", "00101110110011101101010001011010", "00101110000010011101001110001010", "00101101010000011101001010111110", 
			"00101100011101011101000111110110", "00101011101001011101000100110001", "00101010110100111101000001110000", "00101001111111001100111110110010", 
			"00101001001000111100111011111001", "00101000010001101100111001000011", "00100111011001101100110110010001", "00100110100001001100110011100011", 
			"00100101100111101100110000111001", "00100100101101011100101110010011", "00100011110010011100101011110001", "00100010110110111100101001010011", 
			"00100001111010101100100110111001", "00100000111101101100100100100100", "00011111111111111100100010010011", "00011111000001111100100000000110", 
			"00011110000010111100011101111101", "00011101000011101100011011111001", "00011100000011101100011001111010", "00011011000011001100010111111111", 
			"00011010000001111100010110001000", "00011001000000011100010100010110", "00010111111110011100010010101001", "00010110111011111100010001000000", 
			"00010101111000111100001111011100", "00010100110101101100001101111100", "00010011110001101100001100100001", "00010010101101101100001011001011", 
			"00010001101001001100001001111010", "00010000100100001100001000101110", "00001111011110111100000111100110", "00001110011001011100000110100011", 
			"00001101010011101100000101100110", "00001100001101101100000100101101", "00001011000111011100000011111000", "00001010000000111100000011001001", 
			"00001000111010001100000010011111", "00000111110011001100000001111010", "00000110101100001100000001011001", "00000101100100111100000000111110", 
			"00000100011101101100000000100111", "00000011010110011100000000010110", "00000010001110111100000000001001", "00000001000111011100000000000010");
    attribute ram_style: string;
    attribute ram_style of ROM: signal is "block";
begin
    process(clk_a, clk_b)
    begin
        if (rising_edge(clk_a)) then
            if (en_a = '1') then
                data_a_o <= ROM(to_integer(unsigned(addr_a)));
            end if;
        end if;
        
        if (rising_edge(clk_b)) then
            if (en_b = '1') then
                data_b_o <= ROM(to_integer(unsigned(addr_b)));
            end if;
        end if;
    end process;
end Behavioral;
